`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ITESO 
// Engineer:  dariomtz
//////////////////////////////////////////////////////////////////////////////////
module top(
        input [3:0] num,
        output [6:0] disp
    );

    display d(.n(num), .d(disp));

                      
endmodule