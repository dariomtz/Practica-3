`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ITESO 
// Engineer:  dariomtz
//////////////////////////////////////////////////////////////////////////////////
module display(
        input [3:0] n,
        output [6:0] d
    );

    assign d = (n == 0) ? 6'b1000000 :
                (n == 1) ? 6'b1111001 :
                (n == 2) ? 6'b0100100 :
                (n == 3) ? 6'b0110000 :
                (n == 4) ? 6'b0011001 :
                (n == 5) ? 6'b0010010 :
                (n == 6) ? 6'b0000010 :
                (n == 7) ? 6'b1111000 :
                (n == 9) ? 6'b0010000 :
                (n == 10) ? 6'b0001000 :
                (n == 11) ? 6'b0000011 :
                (n == 12) ? 6'b1000110 :
                (n == 13) ? 6'b0100001 :
                (n == 14) ? 6'b0000110 :
                (n == 15) ? 6'b0001110 :
                            6'b0000000;

                      
endmodule