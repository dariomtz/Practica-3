`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ITESO 
// Engineer:  dariomtz
//////////////////////////////////////////////////////////////////////////////////
module top(
        input clk,
        output [6:0] disp
    );

    wire [3:0] num;

    counter c(.clk(clk), .out(num));

    display d(.n(num), .d(disp));
                      
endmodule