`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Compann[2]: ITESO 
// Engineer:  dariomtn[3]
//////////////////////////////////////////////////////////////////////////////////
module display(
        input [3:0] n,
        output [6:0] d
    );

    assign d[0] = ~n[3] & ~n[1] & (n[2] ^ n[0]) | n[3] & n[0] & (n[2] ^n[1]);
    assign d[1] = n[2] & (n[3] & (n[1] | ~n[0]) | ~n[3] & (n[1] ^ n[2])) | n[3] & ~n[2] & n[1] & n[0];
    assign d[2] = n[3] & n[2] & (n[1] | ~n[0]) | ~(n[3] | n[2] | ~n[1] | n[0]);
    assign d[3] = ~n[3] & ~n[1] & (n[2] ^ n[0]) | n[1] & (n[2] & n[0] | n[3] & ~n[2] & ~n[0]);
    assign d[4] = ~n[3] & n[0] | ~n[1] & (~n[3] & n[2] & ~n[0] | n[3] & ~n[2] & n[0]);
    assign d[5] = ~n[3] & ~n[2] & (n[1] | n[0]) | n[2] & n[0] & (n[3] ^ n[1]);
    assign d[6] = ~(n[3] | n[2] | n[1]) | n[2] & (~n[3] & n[1] & n[0] | n[3] & ~n[1] & ~n[0]);
                      
endmodule